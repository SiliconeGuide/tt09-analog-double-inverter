magic
tech sky130A
magscale 1 2
timestamp 1755981816
<< pwell >>
rect 2936 -1374 4694 -926
<< viali >>
rect 2961 546 4728 593
rect 2026 490 2194 538
rect 2984 -996 4678 -932
<< metal1 >>
rect 1159 1011 5242 1286
rect 1159 877 5003 1011
rect 5137 877 5242 1011
rect 1159 836 5242 877
rect 1634 374 1818 836
rect 2016 538 2204 836
rect 2896 593 4780 836
rect 2896 546 2961 593
rect 4728 546 4780 593
rect 2896 540 4780 546
rect 2016 490 2026 538
rect 2194 490 2204 538
rect 2016 474 2204 490
rect 2608 430 4774 482
rect 2608 384 2660 430
rect 1634 278 2094 374
rect 2132 262 2660 384
rect 2843 327 2853 392
rect 2908 327 2918 392
rect 3035 327 3045 392
rect 3100 327 3110 392
rect 3227 327 3237 392
rect 3292 327 3302 392
rect 3419 327 3429 392
rect 3484 327 3494 392
rect 3611 327 3621 392
rect 3676 327 3686 392
rect 3803 327 3813 392
rect 3868 327 3878 392
rect 3995 327 4005 392
rect 4060 327 4070 392
rect 4187 327 4197 392
rect 4252 327 4262 392
rect 4379 327 4389 392
rect 4444 327 4454 392
rect 4571 327 4581 392
rect 4636 327 4646 392
rect 4763 327 4773 392
rect 4828 327 4838 392
rect 1616 132 2146 180
rect 2346 156 2660 262
rect 2939 205 2949 278
rect 3007 205 3017 278
rect 3131 205 3141 278
rect 3199 205 3209 278
rect 3323 205 3333 278
rect 3391 205 3401 278
rect 3515 205 3525 278
rect 3583 205 3593 278
rect 3707 205 3717 278
rect 3775 205 3785 278
rect 3899 205 3909 278
rect 3967 205 3977 278
rect 4091 205 4101 278
rect 4159 205 4169 278
rect 4283 205 4293 278
rect 4351 205 4361 278
rect 4475 205 4485 278
rect 4543 205 4553 278
rect 4667 205 4677 278
rect 4735 205 4745 278
rect 1616 -202 1664 132
rect 2346 104 4700 156
rect 1098 -402 1702 -202
rect 1618 -519 1663 -402
rect 2346 -500 2622 104
rect 5548 -408 5554 -144
rect 5818 -408 6176 -144
rect 1618 -564 2140 -519
rect 2346 -558 4778 -500
rect 1616 -624 1814 -622
rect 1616 -766 2102 -624
rect 2346 -630 2667 -558
rect 2346 -632 2642 -630
rect 2142 -695 2642 -632
rect 2776 -657 2786 -592
rect 2841 -657 2851 -592
rect 2968 -657 2978 -592
rect 3033 -657 3043 -592
rect 3160 -657 3170 -592
rect 3225 -657 3235 -592
rect 3352 -657 3362 -592
rect 3417 -657 3427 -592
rect 3544 -657 3554 -592
rect 3609 -657 3619 -592
rect 3736 -657 3746 -592
rect 3801 -657 3811 -592
rect 3928 -657 3938 -592
rect 3993 -657 4003 -592
rect 4120 -657 4130 -592
rect 4185 -657 4195 -592
rect 4312 -657 4322 -592
rect 4377 -657 4387 -592
rect 4504 -657 4514 -592
rect 4569 -657 4579 -592
rect 4696 -657 4706 -592
rect 4761 -657 4771 -592
rect 2142 -732 2667 -695
rect 1616 -1342 1814 -766
rect 2142 -768 2672 -732
rect 2430 -808 2672 -768
rect 2872 -779 2882 -706
rect 2940 -779 2950 -706
rect 3064 -779 3074 -706
rect 3132 -779 3142 -706
rect 3256 -779 3266 -706
rect 3324 -779 3334 -706
rect 3448 -779 3458 -706
rect 3516 -779 3526 -706
rect 3640 -779 3650 -706
rect 3708 -779 3718 -706
rect 3832 -779 3842 -706
rect 3900 -779 3910 -706
rect 4024 -779 4034 -706
rect 4092 -779 4102 -706
rect 4216 -779 4226 -706
rect 4284 -779 4294 -706
rect 4408 -779 4418 -706
rect 4476 -779 4486 -706
rect 4600 -779 4610 -706
rect 4668 -779 4678 -706
rect 2578 -814 2672 -808
rect 2578 -817 2738 -814
rect 2816 -817 2930 -814
rect 3008 -817 3122 -814
rect 3200 -817 3314 -814
rect 3392 -817 3506 -814
rect 3584 -817 3698 -814
rect 3776 -817 3890 -814
rect 3968 -817 4082 -814
rect 4160 -817 4274 -814
rect 4352 -817 4466 -814
rect 4544 -817 4680 -814
rect 2002 -1312 2220 -858
rect 2578 -866 4680 -817
rect 2578 -870 2672 -866
rect 1998 -1336 2220 -1312
rect 1994 -1342 2220 -1336
rect 2936 -932 4694 -926
rect 2936 -996 2984 -932
rect 4678 -996 4694 -932
rect 2936 -1342 4694 -996
rect 1124 -1498 4913 -1342
rect 5069 -1498 5242 -1342
rect 1124 -1746 5242 -1498
<< via1 >>
rect 5003 877 5137 1011
rect 2853 327 2908 392
rect 3045 327 3100 392
rect 3237 327 3292 392
rect 3429 327 3484 392
rect 3621 327 3676 392
rect 3813 327 3868 392
rect 4005 327 4060 392
rect 4197 327 4252 392
rect 4389 327 4444 392
rect 4581 327 4636 392
rect 4773 327 4828 392
rect 2949 205 3007 278
rect 3141 205 3199 278
rect 3333 205 3391 278
rect 3525 205 3583 278
rect 3717 205 3775 278
rect 3909 205 3967 278
rect 4101 205 4159 278
rect 4293 205 4351 278
rect 4485 205 4543 278
rect 4677 205 4735 278
rect 5554 -408 5818 -144
rect 2786 -657 2841 -592
rect 2978 -657 3033 -592
rect 3170 -657 3225 -592
rect 3362 -657 3417 -592
rect 3554 -657 3609 -592
rect 3746 -657 3801 -592
rect 3938 -657 3993 -592
rect 4130 -657 4185 -592
rect 4322 -657 4377 -592
rect 4514 -657 4569 -592
rect 4706 -657 4761 -592
rect 2882 -779 2940 -706
rect 3074 -779 3132 -706
rect 3266 -779 3324 -706
rect 3458 -779 3516 -706
rect 3650 -779 3708 -706
rect 3842 -779 3900 -706
rect 4034 -779 4092 -706
rect 4226 -779 4284 -706
rect 4418 -779 4476 -706
rect 4610 -779 4668 -706
rect 4913 -1498 5069 -1342
<< metal2 >>
rect 4997 877 5003 1011
rect 5137 877 5143 1011
rect 5003 526 5137 877
rect 2852 400 5137 526
rect 2840 392 5137 400
rect 2840 327 2853 392
rect 2908 327 3045 392
rect 3100 327 3237 392
rect 3292 327 3429 392
rect 3484 327 3621 392
rect 3676 327 3813 392
rect 3868 327 4005 392
rect 4060 327 4197 392
rect 4252 327 4389 392
rect 4444 327 4581 392
rect 4636 327 4773 392
rect 4828 327 4844 392
rect 2840 320 4844 327
rect 2853 317 2908 320
rect 3045 317 3100 320
rect 3237 317 3292 320
rect 3429 317 3484 320
rect 3621 317 3676 320
rect 3813 317 3868 320
rect 4005 317 4060 320
rect 4197 317 4252 320
rect 4389 317 4444 320
rect 4581 317 4636 320
rect 4773 317 4828 320
rect 2949 280 3007 288
rect 3141 280 3199 288
rect 3333 280 3391 288
rect 3525 280 3583 288
rect 3717 280 3775 288
rect 3909 280 3967 288
rect 4101 280 4159 288
rect 4293 280 4351 288
rect 4485 280 4543 288
rect 4677 280 4735 288
rect 2840 278 4874 280
rect 2840 205 2949 278
rect 3007 205 3141 278
rect 3199 205 3333 278
rect 3391 205 3525 278
rect 3583 205 3717 278
rect 3775 205 3909 278
rect 3967 205 4101 278
rect 4159 205 4293 278
rect 4351 205 4485 278
rect 4543 205 4677 278
rect 4735 257 4874 278
rect 4735 256 5129 257
rect 4735 205 5276 256
rect 2840 200 5276 205
rect 2850 118 5276 200
rect 4990 -144 5276 118
rect 5554 -144 5818 -138
rect 4990 -408 5554 -144
rect 2780 -488 4804 -476
rect 4990 -488 5276 -408
rect 5554 -414 5818 -408
rect 2780 -584 5276 -488
rect 2773 -592 5276 -584
rect 2773 -657 2786 -592
rect 2841 -657 2978 -592
rect 3033 -657 3170 -592
rect 3225 -657 3362 -592
rect 3417 -657 3554 -592
rect 3609 -657 3746 -592
rect 3801 -657 3938 -592
rect 3993 -657 4130 -592
rect 4185 -657 4322 -592
rect 4377 -657 4514 -592
rect 4569 -657 4706 -592
rect 4761 -618 5276 -592
rect 4761 -627 5129 -618
rect 4761 -638 4804 -627
rect 4761 -657 4777 -638
rect 2773 -664 4777 -657
rect 2786 -667 2841 -664
rect 2978 -667 3033 -664
rect 3170 -667 3225 -664
rect 3362 -667 3417 -664
rect 3554 -667 3609 -664
rect 3746 -667 3801 -664
rect 3938 -667 3993 -664
rect 4130 -667 4185 -664
rect 4322 -667 4377 -664
rect 4514 -667 4569 -664
rect 4706 -667 4761 -664
rect 2882 -704 2940 -696
rect 3074 -704 3132 -696
rect 3266 -704 3324 -696
rect 3458 -704 3516 -696
rect 3650 -704 3708 -696
rect 3842 -704 3900 -696
rect 4034 -704 4092 -696
rect 4226 -704 4284 -696
rect 4418 -704 4476 -696
rect 4610 -704 4668 -696
rect 2773 -706 4777 -704
rect 2773 -779 2882 -706
rect 2940 -779 3074 -706
rect 3132 -779 3266 -706
rect 3324 -779 3458 -706
rect 3516 -779 3650 -706
rect 3708 -779 3842 -706
rect 3900 -779 4034 -706
rect 4092 -779 4226 -706
rect 4284 -779 4418 -706
rect 4476 -779 4610 -706
rect 4668 -709 4777 -706
rect 4668 -779 5069 -709
rect 2773 -784 5069 -779
rect 2784 -844 5069 -784
rect 4719 -865 5069 -844
rect 4913 -1342 5069 -865
rect 4913 -1504 5069 -1498
use sky130_fd_pr__pfet_01v8_8DVCWJ  sky130_fd_pr__pfet_01v8_8DVCWJ_0
timestamp 1755750298
transform 1 0 3841 0 1 297
box -1127 -319 1127 319
use sky130_fd_pr__pfet_01v8_LGS3BL  XM1
timestamp 1755968424
transform 1 0 2113 0 1 288
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_64Z3AY  XM2
timestamp 1755968424
transform 1 0 2121 0 1 -667
box -211 -279 211 279
use sky130_fd_pr__nfet_01v8_YTLFGX  XM4
timestamp 1755750298
transform 1 0 3775 0 1 -686
box -1127 -310 1127 310
<< labels >>
flabel metal1 1284 964 1484 1164 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 1202 -1572 1402 -1372 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 5908 -378 6108 -178 0 FreeSans 256 0 0 0 output
port 3 nsew
flabel metal1 1098 -402 1298 -202 0 FreeSans 256 0 0 0 input
port 2 nsew
flabel metal1 2358 -708 2506 282 0 FreeSans 320 0 0 0 inverted
<< end >>
