magic
tech sky130A
timestamp 1755742311
<< end >>
