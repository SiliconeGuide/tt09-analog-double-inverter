magic
tech sky130A
magscale 1 2
timestamp 1755970193
<< pwell >>
rect 2936 -1374 4694 -926
<< viali >>
rect 2961 546 4728 593
rect 2026 490 2194 538
rect 2984 -996 4678 -932
<< metal1 >>
rect 1159 836 5242 1286
rect 1634 374 1818 836
rect 2016 538 2204 836
rect 2896 593 4780 836
rect 2896 546 2961 593
rect 4728 546 4780 593
rect 2896 540 4780 546
rect 2016 490 2026 538
rect 2194 490 2204 538
rect 2016 474 2204 490
rect 2608 430 4774 482
rect 2608 384 2660 430
rect 1634 278 2094 374
rect 2132 262 2660 384
rect 1616 132 2146 180
rect 2608 156 2660 262
rect 1616 -202 1664 132
rect 2608 104 4700 156
rect 1098 -402 1702 -202
rect 5908 -378 5944 -178
rect 1618 -519 1663 -402
rect 1618 -564 2140 -519
rect 2609 -558 4778 -500
rect 1616 -624 1814 -622
rect 1616 -766 2102 -624
rect 2609 -632 2667 -558
rect 2142 -732 2667 -632
rect 1616 -1342 1814 -766
rect 2142 -768 2672 -732
rect 2430 -808 2672 -768
rect 2578 -814 2672 -808
rect 2002 -1312 2220 -858
rect 2578 -866 4680 -814
rect 2578 -870 2672 -866
rect 1998 -1336 2220 -1312
rect 1994 -1342 2220 -1336
rect 2936 -932 4694 -926
rect 2936 -996 2984 -932
rect 4678 -996 4694 -932
rect 2936 -1342 4694 -996
rect 1124 -1746 5242 -1342
<< metal2 >>
rect 2840 320 4840 400
rect 2840 200 4840 280
use sky130_fd_pr__pfet_01v8_LGS3BL  XM1
timestamp 1755968424
transform 1 0 2113 0 1 288
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_64Z3AY  XM2
timestamp 1755968424
transform 1 0 2121 0 1 -667
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_8DVCWJ  XM3
timestamp 1755750298
transform 1 0 3841 0 1 297
box -1127 -319 1127 319
use sky130_fd_pr__nfet_01v8_YTLFGX  XM4
timestamp 1755750298
transform 1 0 3775 0 1 -686
box -1127 -310 1127 310
<< labels >>
flabel metal1 1284 964 1484 1164 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 1202 -1572 1402 -1372 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 1098 -402 1298 -202 0 FreeSans 256 0 0 0 input
port 2 nsew
flabel space 5908 -378 6108 -178 0 FreeSans 256 0 0 0 output
port 3 nsew
<< end >>
